`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:54:34 10/17/2019 
// Design Name: 
// Module Name:    alu 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module alu(
	input [31:0] A, 
	input [31:0] B, 
	input [2:0] ALUOp, 
	output [31:0] C
    );

wire [31:0] as_result;

assign C = 
	(ALUOp == 0) ? $unsigned(A) + $unsigned(B) : 
	(ALUOp == 1) ? $unsigned(A) - $unsigned(B) : 
	(ALUOp == 2) ? A & B : 
	(ALUOp == 3) ? A | B : 
	(ALUOp == 4) ? $unsigned(A) >> B : 
	(ALUOp == 5) ? as_result : 
	32'b0;

assign as_result =
        (B[4:0] == 0) ? {{0{A[31]}}, A[31:0]} :
        (B[4:0] == 1) ? {{1{A[31]}}, A[31:1]} :
        (B[4:0] == 2) ? {{2{A[31]}}, A[31:2]} :
        (B[4:0] == 3) ? {{3{A[31]}}, A[31:3]} :
        (B[4:0] == 4) ? {{4{A[31]}}, A[31:4]} :
        (B[4:0] == 5) ? {{5{A[31]}}, A[31:5]} :
        (B[4:0] == 6) ? {{6{A[31]}}, A[31:6]} :
        (B[4:0] == 7) ? {{7{A[31]}}, A[31:7]} :
        (B[4:0] == 8) ? {{8{A[31]}}, A[31:8]} :
        (B[4:0] == 9) ? {{9{A[31]}}, A[31:9]} :
        (B[4:0] == 10) ? {{10{A[31]}}, A[31:10]} :
        (B[4:0] == 11) ? {{11{A[31]}}, A[31:11]} :
        (B[4:0] == 12) ? {{12{A[31]}}, A[31:12]} :
        (B[4:0] == 13) ? {{13{A[31]}}, A[31:13]} :
        (B[4:0] == 14) ? {{14{A[31]}}, A[31:14]} :
        (B[4:0] == 15) ? {{15{A[31]}}, A[31:15]} :
        (B[4:0] == 16) ? {{16{A[31]}}, A[31:16]} :
        (B[4:0] == 17) ? {{17{A[31]}}, A[31:17]} :
        (B[4:0] == 18) ? {{18{A[31]}}, A[31:18]} :
        (B[4:0] == 19) ? {{19{A[31]}}, A[31:19]} :
        (B[4:0] == 20) ? {{20{A[31]}}, A[31:20]} :
        (B[4:0] == 21) ? {{21{A[31]}}, A[31:21]} :
        (B[4:0] == 22) ? {{22{A[31]}}, A[31:22]} :
        (B[4:0] == 23) ? {{23{A[31]}}, A[31:23]} :
        (B[4:0] == 24) ? {{24{A[31]}}, A[31:24]} :
        (B[4:0] == 25) ? {{25{A[31]}}, A[31:25]} :
        (B[4:0] == 26) ? {{26{A[31]}}, A[31:26]} :
        (B[4:0] == 27) ? {{27{A[31]}}, A[31:27]} :
        (B[4:0] == 28) ? {{28{A[31]}}, A[31:28]} :
        (B[4:0] == 29) ? {{29{A[31]}}, A[31:29]} :
        (B[4:0] == 30) ? {{30{A[31]}}, A[31:30]} :
        (B[4:0] == 31) ? {{31{A[31]}}, A[31:31]} :
        {32{A[31]}};

endmodule
