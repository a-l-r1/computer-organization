`include "alu.h"

module alu_tb(
);

initial begin
	$display("hello world");
end

endmodule

