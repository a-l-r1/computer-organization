`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:21:24 09/09/2019 
// Design Name: 
// Module Name:    multi_wire_or_reg_multiple_choice 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module multi_wire_or_reg_multiple_choice(
	input [3:0] a, 
	input [4:7] b, 
	input [8:11] c, 
	output reg [3:0] o1, 
	output reg [4:7] o2
    );

// assign o1[3:0] = a[3:0];
// assign o1[3:0] = b[7:4];
// assign o1[3:0] = b[4:7];
// assign o2[4:7] = c[8:11];
// assign o2[4:7] = c[11:8];

endmodule
