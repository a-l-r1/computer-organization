module cpu(
	input clk
)

/* Control */

control control(
	.clk(clk), 
	.curr_instr()
)

endmodule

